library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity one_pulse_tb is
end entity;

architecture one_pulse_tb_arch of one_pulse_tb is
    begin
end architecture;
