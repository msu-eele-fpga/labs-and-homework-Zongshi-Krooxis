library ieee;
use ieee.std_logic_1164.all;

entity vending_machine_tb is
end entity;


architecture vending_machine_tb_arch of vending_machine_tb is
    begin
end architecture;
