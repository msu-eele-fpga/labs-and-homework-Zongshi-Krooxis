entity timed_counter_tb is
end entity timed_counter_tb;


architecture timed_counter_tb_arch of timed_counter_tb is
    begin
end architecture timed_counter_tb_arch;